
// y(t) = sin(2*pi*F*t), F=261.63Hz, Fs=48000Hz, 16-bit

module lut_C
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 182;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000001000110;
        2: y = 16'b0000000010001101;
        3: y = 16'b0000000011010011;
        4: y = 16'b0000000100011000;
        5: y = 16'b0000000101011110;
        6: y = 16'b0000000110100011;
        7: y = 16'b0000000111100111;
        8: y = 16'b0000001000101011;
        9: y = 16'b0000001001101111;
        10: y = 16'b0000001010110001;
        11: y = 16'b0000001011110011;
        12: y = 16'b0000001100110100;
        13: y = 16'b0000001101110100;
        14: y = 16'b0000001110110011;
        15: y = 16'b0000001111110001;
        16: y = 16'b0000010000101101;
        17: y = 16'b0000010001101001;
        18: y = 16'b0000010010100011;
        19: y = 16'b0000010011011011;
        20: y = 16'b0000010100010010;
        21: y = 16'b0000010101001000;
        22: y = 16'b0000010101111100;
        23: y = 16'b0000010110101110;
        24: y = 16'b0000010111011111;
        25: y = 16'b0000011000001110;
        26: y = 16'b0000011000111011;
        27: y = 16'b0000011001100110;
        28: y = 16'b0000011010001111;
        29: y = 16'b0000011010110111;
        30: y = 16'b0000011011011100;
        31: y = 16'b0000011011111111;
        32: y = 16'b0000011100100000;
        33: y = 16'b0000011100111111;
        34: y = 16'b0000011101011100;
        35: y = 16'b0000011101110110;
        36: y = 16'b0000011110001110;
        37: y = 16'b0000011110100100;
        38: y = 16'b0000011110111000;
        39: y = 16'b0000011111001001;
        40: y = 16'b0000011111011000;
        41: y = 16'b0000011111100101;
        42: y = 16'b0000011111101111;
        43: y = 16'b0000011111110111;
        44: y = 16'b0000011111111100;
        45: y = 16'b0000011111111111;
        46: y = 16'b0000100000000000;
        47: y = 16'b0000011111111110;
        48: y = 16'b0000011111111010;
        49: y = 16'b0000011111110011;
        50: y = 16'b0000011111101010;
        51: y = 16'b0000011111011111;
        52: y = 16'b0000011111010001;
        53: y = 16'b0000011111000001;
        54: y = 16'b0000011110101110;
        55: y = 16'b0000011110011010;
        56: y = 16'b0000011110000010;
        57: y = 16'b0000011101101001;
        58: y = 16'b0000011101001101;
        59: y = 16'b0000011100110000;
        60: y = 16'b0000011100010000;
        61: y = 16'b0000011011101110;
        62: y = 16'b0000011011001001;
        63: y = 16'b0000011010100011;
        64: y = 16'b0000011001111011;
        65: y = 16'b0000011001010001;
        66: y = 16'b0000011000100101;
        67: y = 16'b0000010111110111;
        68: y = 16'b0000010111000111;
        69: y = 16'b0000010110010101;
        70: y = 16'b0000010101100010;
        71: y = 16'b0000010100101101;
        72: y = 16'b0000010011110111;
        73: y = 16'b0000010010111111;
        74: y = 16'b0000010010000110;
        75: y = 16'b0000010001001011;
        76: y = 16'b0000010000001111;
        77: y = 16'b0000001111010010;
        78: y = 16'b0000001110010100;
        79: y = 16'b0000001101010100;
        80: y = 16'b0000001100010100;
        81: y = 16'b0000001011010010;
        82: y = 16'b0000001010010000;
        83: y = 16'b0000001001001101;
        84: y = 16'b0000001000001010;
        85: y = 16'b0000000111000101;
        86: y = 16'b0000000110000000;
        87: y = 16'b0000000100111011;
        88: y = 16'b0000000011110110;
        89: y = 16'b0000000010110000;
        90: y = 16'b0000000001101001;
        91: y = 16'b0000000000100011;
        92: y = 16'b1111111111011101;
        93: y = 16'b1111111110010111;
        94: y = 16'b1111111101010000;
        95: y = 16'b1111111100001010;
        96: y = 16'b1111111011000101;
        97: y = 16'b1111111010000000;
        98: y = 16'b1111111000111011;
        99: y = 16'b1111110111110110;
        100: y = 16'b1111110110110011;
        101: y = 16'b1111110101110000;
        102: y = 16'b1111110100101110;
        103: y = 16'b1111110011101100;
        104: y = 16'b1111110010101100;
        105: y = 16'b1111110001101100;
        106: y = 16'b1111110000101110;
        107: y = 16'b1111101111110001;
        108: y = 16'b1111101110110101;
        109: y = 16'b1111101101111010;
        110: y = 16'b1111101101000001;
        111: y = 16'b1111101100001001;
        112: y = 16'b1111101011010011;
        113: y = 16'b1111101010011110;
        114: y = 16'b1111101001101011;
        115: y = 16'b1111101000111001;
        116: y = 16'b1111101000001001;
        117: y = 16'b1111100111011011;
        118: y = 16'b1111100110101111;
        119: y = 16'b1111100110000101;
        120: y = 16'b1111100101011101;
        121: y = 16'b1111100100110111;
        122: y = 16'b1111100100010010;
        123: y = 16'b1111100011110000;
        124: y = 16'b1111100011010000;
        125: y = 16'b1111100010110011;
        126: y = 16'b1111100010010111;
        127: y = 16'b1111100001111110;
        128: y = 16'b1111100001100110;
        129: y = 16'b1111100001010010;
        130: y = 16'b1111100000111111;
        131: y = 16'b1111100000101111;
        132: y = 16'b1111100000100001;
        133: y = 16'b1111100000010110;
        134: y = 16'b1111100000001101;
        135: y = 16'b1111100000000110;
        136: y = 16'b1111100000000010;
        137: y = 16'b1111100000000000;
        138: y = 16'b1111100000000001;
        139: y = 16'b1111100000000100;
        140: y = 16'b1111100000001001;
        141: y = 16'b1111100000010001;
        142: y = 16'b1111100000011011;
        143: y = 16'b1111100000101000;
        144: y = 16'b1111100000110111;
        145: y = 16'b1111100001001000;
        146: y = 16'b1111100001011100;
        147: y = 16'b1111100001110010;
        148: y = 16'b1111100010001010;
        149: y = 16'b1111100010100100;
        150: y = 16'b1111100011000001;
        151: y = 16'b1111100011100000;
        152: y = 16'b1111100100000001;
        153: y = 16'b1111100100100100;
        154: y = 16'b1111100101001001;
        155: y = 16'b1111100101110001;
        156: y = 16'b1111100110011010;
        157: y = 16'b1111100111000101;
        158: y = 16'b1111100111110010;
        159: y = 16'b1111101000100001;
        160: y = 16'b1111101001010010;
        161: y = 16'b1111101010000100;
        162: y = 16'b1111101010111000;
        163: y = 16'b1111101011101110;
        164: y = 16'b1111101100100101;
        165: y = 16'b1111101101011101;
        166: y = 16'b1111101110010111;
        167: y = 16'b1111101111010011;
        168: y = 16'b1111110000001111;
        169: y = 16'b1111110001001101;
        170: y = 16'b1111110010001100;
        171: y = 16'b1111110011001100;
        172: y = 16'b1111110100001101;
        173: y = 16'b1111110101001111;
        174: y = 16'b1111110110010001;
        175: y = 16'b1111110111010101;
        176: y = 16'b1111111000011001;
        177: y = 16'b1111111001011101;
        178: y = 16'b1111111010100010;
        179: y = 16'b1111111011101000;
        180: y = 16'b1111111100101101;
        181: y = 16'b1111111101110011;
        182: y = 16'b1111111110111010;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=277.18Hz, Fs=48000Hz, 16-bit

module lut_Cs
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 172;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000001001010;
        2: y = 16'b0000000010010101;
        3: y = 16'b0000000011011111;
        4: y = 16'b0000000100101000;
        5: y = 16'b0000000101110010;
        6: y = 16'b0000000110111011;
        7: y = 16'b0000001000000011;
        8: y = 16'b0000001001001011;
        9: y = 16'b0000001010010010;
        10: y = 16'b0000001011011000;
        11: y = 16'b0000001100011101;
        12: y = 16'b0000001101100001;
        13: y = 16'b0000001110100011;
        14: y = 16'b0000001111100101;
        15: y = 16'b0000010000100101;
        16: y = 16'b0000010001100100;
        17: y = 16'b0000010010100010;
        18: y = 16'b0000010011011101;
        19: y = 16'b0000010100011000;
        20: y = 16'b0000010101010000;
        21: y = 16'b0000010110000111;
        22: y = 16'b0000010110111100;
        23: y = 16'b0000010111101111;
        24: y = 16'b0000011000011111;
        25: y = 16'b0000011001001110;
        26: y = 16'b0000011001111011;
        27: y = 16'b0000011010100110;
        28: y = 16'b0000011011001110;
        29: y = 16'b0000011011110100;
        30: y = 16'b0000011100010111;
        31: y = 16'b0000011100111001;
        32: y = 16'b0000011101010111;
        33: y = 16'b0000011101110100;
        34: y = 16'b0000011110001101;
        35: y = 16'b0000011110100101;
        36: y = 16'b0000011110111001;
        37: y = 16'b0000011111001011;
        38: y = 16'b0000011111011011;
        39: y = 16'b0000011111101000;
        40: y = 16'b0000011111110010;
        41: y = 16'b0000011111111001;
        42: y = 16'b0000011111111110;
        43: y = 16'b0000100000000000;
        44: y = 16'b0000011111111111;
        45: y = 16'b0000011111111100;
        46: y = 16'b0000011111110110;
        47: y = 16'b0000011111101101;
        48: y = 16'b0000011111100010;
        49: y = 16'b0000011111010011;
        50: y = 16'b0000011111000011;
        51: y = 16'b0000011110101111;
        52: y = 16'b0000011110011001;
        53: y = 16'b0000011110000001;
        54: y = 16'b0000011101100110;
        55: y = 16'b0000011101001000;
        56: y = 16'b0000011100101000;
        57: y = 16'b0000011100000110;
        58: y = 16'b0000011011100001;
        59: y = 16'b0000011010111010;
        60: y = 16'b0000011010010001;
        61: y = 16'b0000011001100101;
        62: y = 16'b0000011000110111;
        63: y = 16'b0000011000000111;
        64: y = 16'b0000010111010101;
        65: y = 16'b0000010110100010;
        66: y = 16'b0000010101101100;
        67: y = 16'b0000010100110100;
        68: y = 16'b0000010011111011;
        69: y = 16'b0000010011000000;
        70: y = 16'b0000010010000011;
        71: y = 16'b0000010001000101;
        72: y = 16'b0000010000000101;
        73: y = 16'b0000001111000100;
        74: y = 16'b0000001110000010;
        75: y = 16'b0000001100111111;
        76: y = 16'b0000001011111010;
        77: y = 16'b0000001010110101;
        78: y = 16'b0000001001101110;
        79: y = 16'b0000001000100111;
        80: y = 16'b0000000111011111;
        81: y = 16'b0000000110010110;
        82: y = 16'b0000000101001101;
        83: y = 16'b0000000100000100;
        84: y = 16'b0000000010111010;
        85: y = 16'b0000000001110000;
        86: y = 16'b0000000000100101;
        87: y = 16'b1111111111011011;
        88: y = 16'b1111111110010000;
        89: y = 16'b1111111101000110;
        90: y = 16'b1111111011111100;
        91: y = 16'b1111111010110011;
        92: y = 16'b1111111001101010;
        93: y = 16'b1111111000100001;
        94: y = 16'b1111110111011001;
        95: y = 16'b1111110110010010;
        96: y = 16'b1111110101001011;
        97: y = 16'b1111110100000110;
        98: y = 16'b1111110011000001;
        99: y = 16'b1111110001111110;
        100: y = 16'b1111110000111100;
        101: y = 16'b1111101111111011;
        102: y = 16'b1111101110111011;
        103: y = 16'b1111101101111101;
        104: y = 16'b1111101101000000;
        105: y = 16'b1111101100000101;
        106: y = 16'b1111101011001100;
        107: y = 16'b1111101010010100;
        108: y = 16'b1111101001011110;
        109: y = 16'b1111101000101011;
        110: y = 16'b1111100111111001;
        111: y = 16'b1111100111001001;
        112: y = 16'b1111100110011011;
        113: y = 16'b1111100101101111;
        114: y = 16'b1111100101000110;
        115: y = 16'b1111100100011111;
        116: y = 16'b1111100011111010;
        117: y = 16'b1111100011011000;
        118: y = 16'b1111100010111000;
        119: y = 16'b1111100010011010;
        120: y = 16'b1111100001111111;
        121: y = 16'b1111100001100111;
        122: y = 16'b1111100001010001;
        123: y = 16'b1111100000111101;
        124: y = 16'b1111100000101101;
        125: y = 16'b1111100000011110;
        126: y = 16'b1111100000010011;
        127: y = 16'b1111100000001010;
        128: y = 16'b1111100000000100;
        129: y = 16'b1111100000000001;
        130: y = 16'b1111100000000000;
        131: y = 16'b1111100000000010;
        132: y = 16'b1111100000000111;
        133: y = 16'b1111100000001110;
        134: y = 16'b1111100000011000;
        135: y = 16'b1111100000100101;
        136: y = 16'b1111100000110101;
        137: y = 16'b1111100001000111;
        138: y = 16'b1111100001011011;
        139: y = 16'b1111100001110011;
        140: y = 16'b1111100010001100;
        141: y = 16'b1111100010101001;
        142: y = 16'b1111100011000111;
        143: y = 16'b1111100011101001;
        144: y = 16'b1111100100001100;
        145: y = 16'b1111100100110010;
        146: y = 16'b1111100101011010;
        147: y = 16'b1111100110000101;
        148: y = 16'b1111100110110010;
        149: y = 16'b1111100111100001;
        150: y = 16'b1111101000010001;
        151: y = 16'b1111101001000100;
        152: y = 16'b1111101001111001;
        153: y = 16'b1111101010110000;
        154: y = 16'b1111101011101000;
        155: y = 16'b1111101100100011;
        156: y = 16'b1111101101011110;
        157: y = 16'b1111101110011100;
        158: y = 16'b1111101111011011;
        159: y = 16'b1111110000011011;
        160: y = 16'b1111110001011101;
        161: y = 16'b1111110010011111;
        162: y = 16'b1111110011100011;
        163: y = 16'b1111110100101000;
        164: y = 16'b1111110101101110;
        165: y = 16'b1111110110110101;
        166: y = 16'b1111110111111101;
        167: y = 16'b1111111001000101;
        168: y = 16'b1111111010001110;
        169: y = 16'b1111111011011000;
        170: y = 16'b1111111100100001;
        171: y = 16'b1111111101101011;
        172: y = 16'b1111111110110110;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=293.66Hz, Fs=48000Hz, 16-bit

module lut_D
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 162;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000001001111;
        2: y = 16'b0000000010011110;
        3: y = 16'b0000000011101100;
        4: y = 16'b0000000100111011;
        5: y = 16'b0000000110001000;
        6: y = 16'b0000000111010101;
        7: y = 16'b0000001000100010;
        8: y = 16'b0000001001101110;
        9: y = 16'b0000001010111000;
        10: y = 16'b0000001100000010;
        11: y = 16'b0000001101001011;
        12: y = 16'b0000001110010010;
        13: y = 16'b0000001111011000;
        14: y = 16'b0000010000011100;
        15: y = 16'b0000010001011111;
        16: y = 16'b0000010010100001;
        17: y = 16'b0000010011100000;
        18: y = 16'b0000010100011110;
        19: y = 16'b0000010101011001;
        20: y = 16'b0000010110010011;
        21: y = 16'b0000010111001011;
        22: y = 16'b0000011000000000;
        23: y = 16'b0000011000110011;
        24: y = 16'b0000011001100100;
        25: y = 16'b0000011010010010;
        26: y = 16'b0000011010111110;
        27: y = 16'b0000011011100111;
        28: y = 16'b0000011100001110;
        29: y = 16'b0000011100110001;
        30: y = 16'b0000011101010011;
        31: y = 16'b0000011101110001;
        32: y = 16'b0000011110001101;
        33: y = 16'b0000011110100101;
        34: y = 16'b0000011110111011;
        35: y = 16'b0000011111001110;
        36: y = 16'b0000011111011110;
        37: y = 16'b0000011111101011;
        38: y = 16'b0000011111110100;
        39: y = 16'b0000011111111011;
        40: y = 16'b0000011111111111;
        41: y = 16'b0000100000000000;
        42: y = 16'b0000011111111110;
        43: y = 16'b0000011111111000;
        44: y = 16'b0000011111110000;
        45: y = 16'b0000011111100101;
        46: y = 16'b0000011111010110;
        47: y = 16'b0000011111000101;
        48: y = 16'b0000011110110000;
        49: y = 16'b0000011110011001;
        50: y = 16'b0000011101111111;
        51: y = 16'b0000011101100010;
        52: y = 16'b0000011101000010;
        53: y = 16'b0000011100100000;
        54: y = 16'b0000011011111011;
        55: y = 16'b0000011011010011;
        56: y = 16'b0000011010101000;
        57: y = 16'b0000011001111011;
        58: y = 16'b0000011001001100;
        59: y = 16'b0000011000011010;
        60: y = 16'b0000010111100110;
        61: y = 16'b0000010110101111;
        62: y = 16'b0000010101110110;
        63: y = 16'b0000010100111100;
        64: y = 16'b0000010011111111;
        65: y = 16'b0000010011000000;
        66: y = 16'b0000010010000000;
        67: y = 16'b0000010000111110;
        68: y = 16'b0000001111111010;
        69: y = 16'b0000001110110101;
        70: y = 16'b0000001101101110;
        71: y = 16'b0000001100100110;
        72: y = 16'b0000001011011101;
        73: y = 16'b0000001010010011;
        74: y = 16'b0000001001001000;
        75: y = 16'b0000000111111100;
        76: y = 16'b0000000110101111;
        77: y = 16'b0000000101100001;
        78: y = 16'b0000000100010011;
        79: y = 16'b0000000011000101;
        80: y = 16'b0000000001110110;
        81: y = 16'b0000000000100111;
        82: y = 16'b1111111111011001;
        83: y = 16'b1111111110001010;
        84: y = 16'b1111111100111011;
        85: y = 16'b1111111011101101;
        86: y = 16'b1111111010011111;
        87: y = 16'b1111111001010001;
        88: y = 16'b1111111000000100;
        89: y = 16'b1111110110111000;
        90: y = 16'b1111110101101101;
        91: y = 16'b1111110100100011;
        92: y = 16'b1111110011011010;
        93: y = 16'b1111110010010010;
        94: y = 16'b1111110001001011;
        95: y = 16'b1111110000000110;
        96: y = 16'b1111101111000010;
        97: y = 16'b1111101110000000;
        98: y = 16'b1111101101000000;
        99: y = 16'b1111101100000001;
        100: y = 16'b1111101011000100;
        101: y = 16'b1111101010001010;
        102: y = 16'b1111101001010001;
        103: y = 16'b1111101000011010;
        104: y = 16'b1111100111100110;
        105: y = 16'b1111100110110100;
        106: y = 16'b1111100110000101;
        107: y = 16'b1111100101011000;
        108: y = 16'b1111100100101101;
        109: y = 16'b1111100100000101;
        110: y = 16'b1111100011100000;
        111: y = 16'b1111100010111110;
        112: y = 16'b1111100010011110;
        113: y = 16'b1111100010000001;
        114: y = 16'b1111100001100111;
        115: y = 16'b1111100001010000;
        116: y = 16'b1111100000111011;
        117: y = 16'b1111100000101010;
        118: y = 16'b1111100000011011;
        119: y = 16'b1111100000010000;
        120: y = 16'b1111100000001000;
        121: y = 16'b1111100000000010;
        122: y = 16'b1111100000000000;
        123: y = 16'b1111100000000001;
        124: y = 16'b1111100000000101;
        125: y = 16'b1111100000001100;
        126: y = 16'b1111100000010101;
        127: y = 16'b1111100000100010;
        128: y = 16'b1111100000110010;
        129: y = 16'b1111100001000101;
        130: y = 16'b1111100001011011;
        131: y = 16'b1111100001110011;
        132: y = 16'b1111100010001111;
        133: y = 16'b1111100010101101;
        134: y = 16'b1111100011001111;
        135: y = 16'b1111100011110010;
        136: y = 16'b1111100100011001;
        137: y = 16'b1111100101000010;
        138: y = 16'b1111100101101110;
        139: y = 16'b1111100110011100;
        140: y = 16'b1111100111001101;
        141: y = 16'b1111101000000000;
        142: y = 16'b1111101000110101;
        143: y = 16'b1111101001101101;
        144: y = 16'b1111101010100111;
        145: y = 16'b1111101011100010;
        146: y = 16'b1111101100100000;
        147: y = 16'b1111101101011111;
        148: y = 16'b1111101110100001;
        149: y = 16'b1111101111100100;
        150: y = 16'b1111110000101000;
        151: y = 16'b1111110001101110;
        152: y = 16'b1111110010110101;
        153: y = 16'b1111110011111110;
        154: y = 16'b1111110101001000;
        155: y = 16'b1111110110010010;
        156: y = 16'b1111110111011110;
        157: y = 16'b1111111000101011;
        158: y = 16'b1111111001111000;
        159: y = 16'b1111111011000101;
        160: y = 16'b1111111100010100;
        161: y = 16'b1111111101100010;
        162: y = 16'b1111111110110001;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=311.13Hz, Fs=48000Hz, 16-bit

module lut_Ds
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 153;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000001010100;
        2: y = 16'b0000000010100111;
        3: y = 16'b0000000011111010;
        4: y = 16'b0000000101001101;
        5: y = 16'b0000000110011111;
        6: y = 16'b0000000111110000;
        7: y = 16'b0000001001000001;
        8: y = 16'b0000001010010001;
        9: y = 16'b0000001011011111;
        10: y = 16'b0000001100101101;
        11: y = 16'b0000001101111001;
        12: y = 16'b0000001111000011;
        13: y = 16'b0000010000001100;
        14: y = 16'b0000010001010011;
        15: y = 16'b0000010010011001;
        16: y = 16'b0000010011011100;
        17: y = 16'b0000010100011101;
        18: y = 16'b0000010101011100;
        19: y = 16'b0000010110011001;
        20: y = 16'b0000010111010100;
        21: y = 16'b0000011000001100;
        22: y = 16'b0000011001000001;
        23: y = 16'b0000011001110100;
        24: y = 16'b0000011010100100;
        25: y = 16'b0000011011010001;
        26: y = 16'b0000011011111011;
        27: y = 16'b0000011100100011;
        28: y = 16'b0000011101000111;
        29: y = 16'b0000011101101000;
        30: y = 16'b0000011110000110;
        31: y = 16'b0000011110100001;
        32: y = 16'b0000011110111000;
        33: y = 16'b0000011111001101;
        34: y = 16'b0000011111011110;
        35: y = 16'b0000011111101011;
        36: y = 16'b0000011111110101;
        37: y = 16'b0000011111111100;
        38: y = 16'b0000100000000000;
        39: y = 16'b0000100000000000;
        40: y = 16'b0000011111111100;
        41: y = 16'b0000011111110101;
        42: y = 16'b0000011111101011;
        43: y = 16'b0000011111011110;
        44: y = 16'b0000011111001101;
        45: y = 16'b0000011110111000;
        46: y = 16'b0000011110100001;
        47: y = 16'b0000011110000110;
        48: y = 16'b0000011101101000;
        49: y = 16'b0000011101000111;
        50: y = 16'b0000011100100011;
        51: y = 16'b0000011011111011;
        52: y = 16'b0000011011010001;
        53: y = 16'b0000011010100100;
        54: y = 16'b0000011001110100;
        55: y = 16'b0000011001000001;
        56: y = 16'b0000011000001100;
        57: y = 16'b0000010111010100;
        58: y = 16'b0000010110011001;
        59: y = 16'b0000010101011100;
        60: y = 16'b0000010100011101;
        61: y = 16'b0000010011011100;
        62: y = 16'b0000010010011001;
        63: y = 16'b0000010001010011;
        64: y = 16'b0000010000001100;
        65: y = 16'b0000001111000011;
        66: y = 16'b0000001101111001;
        67: y = 16'b0000001100101101;
        68: y = 16'b0000001011011111;
        69: y = 16'b0000001010010001;
        70: y = 16'b0000001001000001;
        71: y = 16'b0000000111110000;
        72: y = 16'b0000000110011111;
        73: y = 16'b0000000101001101;
        74: y = 16'b0000000011111010;
        75: y = 16'b0000000010100111;
        76: y = 16'b0000000001010100;
        77: y = 16'b0000000000000000;
        78: y = 16'b1111111110101100;
        79: y = 16'b1111111101011001;
        80: y = 16'b1111111100000110;
        81: y = 16'b1111111010110011;
        82: y = 16'b1111111001100001;
        83: y = 16'b1111111000010000;
        84: y = 16'b1111110110111111;
        85: y = 16'b1111110101101111;
        86: y = 16'b1111110100100001;
        87: y = 16'b1111110011010011;
        88: y = 16'b1111110010000111;
        89: y = 16'b1111110000111101;
        90: y = 16'b1111101111110100;
        91: y = 16'b1111101110101101;
        92: y = 16'b1111101101100111;
        93: y = 16'b1111101100100100;
        94: y = 16'b1111101011100011;
        95: y = 16'b1111101010100100;
        96: y = 16'b1111101001100111;
        97: y = 16'b1111101000101100;
        98: y = 16'b1111100111110100;
        99: y = 16'b1111100110111111;
        100: y = 16'b1111100110001100;
        101: y = 16'b1111100101011100;
        102: y = 16'b1111100100101111;
        103: y = 16'b1111100100000101;
        104: y = 16'b1111100011011101;
        105: y = 16'b1111100010111001;
        106: y = 16'b1111100010011000;
        107: y = 16'b1111100001111010;
        108: y = 16'b1111100001011111;
        109: y = 16'b1111100001001000;
        110: y = 16'b1111100000110011;
        111: y = 16'b1111100000100010;
        112: y = 16'b1111100000010101;
        113: y = 16'b1111100000001011;
        114: y = 16'b1111100000000100;
        115: y = 16'b1111100000000000;
        116: y = 16'b1111100000000000;
        117: y = 16'b1111100000000100;
        118: y = 16'b1111100000001011;
        119: y = 16'b1111100000010101;
        120: y = 16'b1111100000100010;
        121: y = 16'b1111100000110011;
        122: y = 16'b1111100001001000;
        123: y = 16'b1111100001011111;
        124: y = 16'b1111100001111010;
        125: y = 16'b1111100010011000;
        126: y = 16'b1111100010111001;
        127: y = 16'b1111100011011101;
        128: y = 16'b1111100100000101;
        129: y = 16'b1111100100101111;
        130: y = 16'b1111100101011100;
        131: y = 16'b1111100110001100;
        132: y = 16'b1111100110111111;
        133: y = 16'b1111100111110100;
        134: y = 16'b1111101000101100;
        135: y = 16'b1111101001100111;
        136: y = 16'b1111101010100100;
        137: y = 16'b1111101011100011;
        138: y = 16'b1111101100100100;
        139: y = 16'b1111101101100111;
        140: y = 16'b1111101110101101;
        141: y = 16'b1111101111110100;
        142: y = 16'b1111110000111101;
        143: y = 16'b1111110010000111;
        144: y = 16'b1111110011010011;
        145: y = 16'b1111110100100001;
        146: y = 16'b1111110101101111;
        147: y = 16'b1111110110111111;
        148: y = 16'b1111111000010000;
        149: y = 16'b1111111001100001;
        150: y = 16'b1111111010110011;
        151: y = 16'b1111111100000110;
        152: y = 16'b1111111101011001;
        153: y = 16'b1111111110101100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=329.63Hz, Fs=48000Hz, 16-bit

module lut_E
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 144;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000001011001;
        2: y = 16'b0000000010110001;
        3: y = 16'b0000000100001001;
        4: y = 16'b0000000101100001;
        5: y = 16'b0000000110111000;
        6: y = 16'b0000001000001110;
        7: y = 16'b0000001001100100;
        8: y = 16'b0000001010111000;
        9: y = 16'b0000001100001011;
        10: y = 16'b0000001101011100;
        11: y = 16'b0000001110101100;
        12: y = 16'b0000001111111010;
        13: y = 16'b0000010001000110;
        14: y = 16'b0000010010010000;
        15: y = 16'b0000010011010111;
        16: y = 16'b0000010100011101;
        17: y = 16'b0000010101100000;
        18: y = 16'b0000010110100000;
        19: y = 16'b0000010111011110;
        20: y = 16'b0000011000011001;
        21: y = 16'b0000011001010001;
        22: y = 16'b0000011010000110;
        23: y = 16'b0000011010111000;
        24: y = 16'b0000011011100110;
        25: y = 16'b0000011100010001;
        26: y = 16'b0000011100111001;
        27: y = 16'b0000011101011110;
        28: y = 16'b0000011101111110;
        29: y = 16'b0000011110011100;
        30: y = 16'b0000011110110101;
        31: y = 16'b0000011111001011;
        32: y = 16'b0000011111011101;
        33: y = 16'b0000011111101100;
        34: y = 16'b0000011111110110;
        35: y = 16'b0000011111111101;
        36: y = 16'b0000100000000000;
        37: y = 16'b0000011111111111;
        38: y = 16'b0000011111111010;
        39: y = 16'b0000011111110001;
        40: y = 16'b0000011111100101;
        41: y = 16'b0000011111010101;
        42: y = 16'b0000011111000001;
        43: y = 16'b0000011110101001;
        44: y = 16'b0000011110001110;
        45: y = 16'b0000011101101110;
        46: y = 16'b0000011101001100;
        47: y = 16'b0000011100100110;
        48: y = 16'b0000011011111100;
        49: y = 16'b0000011011001111;
        50: y = 16'b0000011010011111;
        51: y = 16'b0000011001101100;
        52: y = 16'b0000011000110101;
        53: y = 16'b0000010111111100;
        54: y = 16'b0000010110111111;
        55: y = 16'b0000010110000000;
        56: y = 16'b0000010100111111;
        57: y = 16'b0000010011111010;
        58: y = 16'b0000010010110100;
        59: y = 16'b0000010001101011;
        60: y = 16'b0000010000100000;
        61: y = 16'b0000001111010011;
        62: y = 16'b0000001110000100;
        63: y = 16'b0000001100110011;
        64: y = 16'b0000001011100001;
        65: y = 16'b0000001010001110;
        66: y = 16'b0000001000111001;
        67: y = 16'b0000000111100011;
        68: y = 16'b0000000110001101;
        69: y = 16'b0000000100110101;
        70: y = 16'b0000000011011101;
        71: y = 16'b0000000010000101;
        72: y = 16'b0000000000101100;
        73: y = 16'b1111111111010100;
        74: y = 16'b1111111101111011;
        75: y = 16'b1111111100100011;
        76: y = 16'b1111111011001011;
        77: y = 16'b1111111001110011;
        78: y = 16'b1111111000011101;
        79: y = 16'b1111110111000111;
        80: y = 16'b1111110101110010;
        81: y = 16'b1111110100011111;
        82: y = 16'b1111110011001101;
        83: y = 16'b1111110001111100;
        84: y = 16'b1111110000101101;
        85: y = 16'b1111101111100000;
        86: y = 16'b1111101110010101;
        87: y = 16'b1111101101001100;
        88: y = 16'b1111101100000110;
        89: y = 16'b1111101011000001;
        90: y = 16'b1111101010000000;
        91: y = 16'b1111101001000001;
        92: y = 16'b1111101000000100;
        93: y = 16'b1111100111001011;
        94: y = 16'b1111100110010100;
        95: y = 16'b1111100101100001;
        96: y = 16'b1111100100110001;
        97: y = 16'b1111100100000100;
        98: y = 16'b1111100011011010;
        99: y = 16'b1111100010110100;
        100: y = 16'b1111100010010010;
        101: y = 16'b1111100001110010;
        102: y = 16'b1111100001010111;
        103: y = 16'b1111100000111111;
        104: y = 16'b1111100000101011;
        105: y = 16'b1111100000011011;
        106: y = 16'b1111100000001111;
        107: y = 16'b1111100000000110;
        108: y = 16'b1111100000000001;
        109: y = 16'b1111100000000000;
        110: y = 16'b1111100000000011;
        111: y = 16'b1111100000001010;
        112: y = 16'b1111100000010100;
        113: y = 16'b1111100000100011;
        114: y = 16'b1111100000110101;
        115: y = 16'b1111100001001011;
        116: y = 16'b1111100001100100;
        117: y = 16'b1111100010000010;
        118: y = 16'b1111100010100010;
        119: y = 16'b1111100011000111;
        120: y = 16'b1111100011101111;
        121: y = 16'b1111100100011010;
        122: y = 16'b1111100101001000;
        123: y = 16'b1111100101111010;
        124: y = 16'b1111100110101111;
        125: y = 16'b1111100111100111;
        126: y = 16'b1111101000100010;
        127: y = 16'b1111101001100000;
        128: y = 16'b1111101010100000;
        129: y = 16'b1111101011100011;
        130: y = 16'b1111101100101001;
        131: y = 16'b1111101101110000;
        132: y = 16'b1111101110111010;
        133: y = 16'b1111110000000110;
        134: y = 16'b1111110001010100;
        135: y = 16'b1111110010100100;
        136: y = 16'b1111110011110101;
        137: y = 16'b1111110101001000;
        138: y = 16'b1111110110011100;
        139: y = 16'b1111110111110010;
        140: y = 16'b1111111001001000;
        141: y = 16'b1111111010011111;
        142: y = 16'b1111111011110111;
        143: y = 16'b1111111101001111;
        144: y = 16'b1111111110100111;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=349.23Hz, Fs=48000Hz, 16-bit

module lut_F
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 136;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000001011110;
        2: y = 16'b0000000010111100;
        3: y = 16'b0000000100011001;
        4: y = 16'b0000000101110110;
        5: y = 16'b0000000111010010;
        6: y = 16'b0000001000101100;
        7: y = 16'b0000001010000110;
        8: y = 16'b0000001011011111;
        9: y = 16'b0000001100110110;
        10: y = 16'b0000001110001011;
        11: y = 16'b0000001111011110;
        12: y = 16'b0000010000101111;
        13: y = 16'b0000010001111110;
        14: y = 16'b0000010011001010;
        15: y = 16'b0000010100010100;
        16: y = 16'b0000010101011100;
        17: y = 16'b0000010110100000;
        18: y = 16'b0000010111100001;
        19: y = 16'b0000011000011111;
        20: y = 16'b0000011001011010;
        21: y = 16'b0000011010010001;
        22: y = 16'b0000011011000101;
        23: y = 16'b0000011011110101;
        24: y = 16'b0000011100100010;
        25: y = 16'b0000011101001010;
        26: y = 16'b0000011101101111;
        27: y = 16'b0000011110010000;
        28: y = 16'b0000011110101100;
        29: y = 16'b0000011111000101;
        30: y = 16'b0000011111011001;
        31: y = 16'b0000011111101001;
        32: y = 16'b0000011111110101;
        33: y = 16'b0000011111111101;
        34: y = 16'b0000100000000000;
        35: y = 16'b0000011111111111;
        36: y = 16'b0000011111111001;
        37: y = 16'b0000011111110000;
        38: y = 16'b0000011111100010;
        39: y = 16'b0000011111010000;
        40: y = 16'b0000011110111001;
        41: y = 16'b0000011110011111;
        42: y = 16'b0000011110000000;
        43: y = 16'b0000011101011101;
        44: y = 16'b0000011100110111;
        45: y = 16'b0000011100001100;
        46: y = 16'b0000011011011110;
        47: y = 16'b0000011010101100;
        48: y = 16'b0000011001110110;
        49: y = 16'b0000011000111101;
        50: y = 16'b0000011000000000;
        51: y = 16'b0000010111000001;
        52: y = 16'b0000010101111110;
        53: y = 16'b0000010100111000;
        54: y = 16'b0000010011110000;
        55: y = 16'b0000010010100100;
        56: y = 16'b0000010001010111;
        57: y = 16'b0000010000000111;
        58: y = 16'b0000001110110101;
        59: y = 16'b0000001101100000;
        60: y = 16'b0000001100001010;
        61: y = 16'b0000001010110011;
        62: y = 16'b0000001001011010;
        63: y = 16'b0000000111111111;
        64: y = 16'b0000000110100100;
        65: y = 16'b0000000101000111;
        66: y = 16'b0000000011101010;
        67: y = 16'b0000000010001101;
        68: y = 16'b0000000000101111;
        69: y = 16'b1111111111010001;
        70: y = 16'b1111111101110011;
        71: y = 16'b1111111100010110;
        72: y = 16'b1111111010111001;
        73: y = 16'b1111111001011100;
        74: y = 16'b1111111000000001;
        75: y = 16'b1111110110100110;
        76: y = 16'b1111110101001101;
        77: y = 16'b1111110011110110;
        78: y = 16'b1111110010100000;
        79: y = 16'b1111110001001011;
        80: y = 16'b1111101111111001;
        81: y = 16'b1111101110101001;
        82: y = 16'b1111101101011100;
        83: y = 16'b1111101100010000;
        84: y = 16'b1111101011001000;
        85: y = 16'b1111101010000010;
        86: y = 16'b1111101000111111;
        87: y = 16'b1111101000000000;
        88: y = 16'b1111100111000011;
        89: y = 16'b1111100110001010;
        90: y = 16'b1111100101010100;
        91: y = 16'b1111100100100010;
        92: y = 16'b1111100011110100;
        93: y = 16'b1111100011001001;
        94: y = 16'b1111100010100011;
        95: y = 16'b1111100010000000;
        96: y = 16'b1111100001100001;
        97: y = 16'b1111100001000111;
        98: y = 16'b1111100000110000;
        99: y = 16'b1111100000011110;
        100: y = 16'b1111100000010000;
        101: y = 16'b1111100000000111;
        102: y = 16'b1111100000000001;
        103: y = 16'b1111100000000000;
        104: y = 16'b1111100000000011;
        105: y = 16'b1111100000001011;
        106: y = 16'b1111100000010111;
        107: y = 16'b1111100000100111;
        108: y = 16'b1111100000111011;
        109: y = 16'b1111100001010100;
        110: y = 16'b1111100001110000;
        111: y = 16'b1111100010010001;
        112: y = 16'b1111100010110110;
        113: y = 16'b1111100011011110;
        114: y = 16'b1111100100001011;
        115: y = 16'b1111100100111011;
        116: y = 16'b1111100101101111;
        117: y = 16'b1111100110100110;
        118: y = 16'b1111100111100001;
        119: y = 16'b1111101000011111;
        120: y = 16'b1111101001100000;
        121: y = 16'b1111101010100100;
        122: y = 16'b1111101011101100;
        123: y = 16'b1111101100110110;
        124: y = 16'b1111101110000010;
        125: y = 16'b1111101111010001;
        126: y = 16'b1111110000100010;
        127: y = 16'b1111110001110101;
        128: y = 16'b1111110011001010;
        129: y = 16'b1111110100100001;
        130: y = 16'b1111110101111010;
        131: y = 16'b1111110111010100;
        132: y = 16'b1111111000101110;
        133: y = 16'b1111111010001010;
        134: y = 16'b1111111011100111;
        135: y = 16'b1111111101000100;
        136: y = 16'b1111111110100010;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=369.99Hz, Fs=48000Hz, 16-bit

module lut_Fs
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 128;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000001100100;
        2: y = 16'b0000000011000111;
        3: y = 16'b0000000100101010;
        4: y = 16'b0000000110001100;
        5: y = 16'b0000000111101110;
        6: y = 16'b0000001001001110;
        7: y = 16'b0000001010101101;
        8: y = 16'b0000001100001010;
        9: y = 16'b0000001101100101;
        10: y = 16'b0000001110111111;
        11: y = 16'b0000010000010101;
        12: y = 16'b0000010001101010;
        13: y = 16'b0000010010111100;
        14: y = 16'b0000010100001011;
        15: y = 16'b0000010101010111;
        16: y = 16'b0000010110011111;
        17: y = 16'b0000010111100100;
        18: y = 16'b0000011000100110;
        19: y = 16'b0000011001100100;
        20: y = 16'b0000011010011110;
        21: y = 16'b0000011011010100;
        22: y = 16'b0000011100000110;
        23: y = 16'b0000011100110100;
        24: y = 16'b0000011101011101;
        25: y = 16'b0000011110000010;
        26: y = 16'b0000011110100010;
        27: y = 16'b0000011110111101;
        28: y = 16'b0000011111010100;
        29: y = 16'b0000011111100110;
        30: y = 16'b0000011111110100;
        31: y = 16'b0000011111111100;
        32: y = 16'b0000100000000000;
        33: y = 16'b0000011111111111;
        34: y = 16'b0000011111111001;
        35: y = 16'b0000011111101110;
        36: y = 16'b0000011111011110;
        37: y = 16'b0000011111001001;
        38: y = 16'b0000011110110000;
        39: y = 16'b0000011110010010;
        40: y = 16'b0000011101110000;
        41: y = 16'b0000011101001001;
        42: y = 16'b0000011100011101;
        43: y = 16'b0000011011101110;
        44: y = 16'b0000011010111010;
        45: y = 16'b0000011010000010;
        46: y = 16'b0000011001000110;
        47: y = 16'b0000011000000110;
        48: y = 16'b0000010111000010;
        49: y = 16'b0000010101111011;
        50: y = 16'b0000010100110001;
        51: y = 16'b0000010011100100;
        52: y = 16'b0000010010010011;
        53: y = 16'b0000010001000000;
        54: y = 16'b0000001111101010;
        55: y = 16'b0000001110010010;
        56: y = 16'b0000001100111000;
        57: y = 16'b0000001011011100;
        58: y = 16'b0000001001111110;
        59: y = 16'b0000001000011110;
        60: y = 16'b0000000110111101;
        61: y = 16'b0000000101011011;
        62: y = 16'b0000000011111001;
        63: y = 16'b0000000010010101;
        64: y = 16'b0000000000110010;
        65: y = 16'b1111111111001110;
        66: y = 16'b1111111101101011;
        67: y = 16'b1111111100000111;
        68: y = 16'b1111111010100101;
        69: y = 16'b1111111001000011;
        70: y = 16'b1111110111100010;
        71: y = 16'b1111110110000010;
        72: y = 16'b1111110100100100;
        73: y = 16'b1111110011001000;
        74: y = 16'b1111110001101110;
        75: y = 16'b1111110000010110;
        76: y = 16'b1111101111000000;
        77: y = 16'b1111101101101101;
        78: y = 16'b1111101100011100;
        79: y = 16'b1111101011001111;
        80: y = 16'b1111101010000101;
        81: y = 16'b1111101000111110;
        82: y = 16'b1111100111111010;
        83: y = 16'b1111100110111010;
        84: y = 16'b1111100101111110;
        85: y = 16'b1111100101000110;
        86: y = 16'b1111100100010010;
        87: y = 16'b1111100011100011;
        88: y = 16'b1111100010110111;
        89: y = 16'b1111100010010000;
        90: y = 16'b1111100001101110;
        91: y = 16'b1111100001010000;
        92: y = 16'b1111100000110111;
        93: y = 16'b1111100000100010;
        94: y = 16'b1111100000010010;
        95: y = 16'b1111100000000111;
        96: y = 16'b1111100000000001;
        97: y = 16'b1111100000000000;
        98: y = 16'b1111100000000100;
        99: y = 16'b1111100000001100;
        100: y = 16'b1111100000011010;
        101: y = 16'b1111100000101100;
        102: y = 16'b1111100001000011;
        103: y = 16'b1111100001011110;
        104: y = 16'b1111100001111110;
        105: y = 16'b1111100010100011;
        106: y = 16'b1111100011001100;
        107: y = 16'b1111100011111010;
        108: y = 16'b1111100100101100;
        109: y = 16'b1111100101100010;
        110: y = 16'b1111100110011100;
        111: y = 16'b1111100111011010;
        112: y = 16'b1111101000011100;
        113: y = 16'b1111101001100001;
        114: y = 16'b1111101010101001;
        115: y = 16'b1111101011110101;
        116: y = 16'b1111101101000100;
        117: y = 16'b1111101110010110;
        118: y = 16'b1111101111101011;
        119: y = 16'b1111110001000001;
        120: y = 16'b1111110010011011;
        121: y = 16'b1111110011110110;
        122: y = 16'b1111110101010011;
        123: y = 16'b1111110110110010;
        124: y = 16'b1111111000010010;
        125: y = 16'b1111111001110100;
        126: y = 16'b1111111011010110;
        127: y = 16'b1111111100111001;
        128: y = 16'b1111111110011100;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=392.0Hz, Fs=48000Hz, 16-bit

module lut_G
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 121;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000001101001;
        2: y = 16'b0000000011010011;
        3: y = 16'b0000000100111011;
        4: y = 16'b0000000110100011;
        5: y = 16'b0000001000001010;
        6: y = 16'b0000001001101111;
        7: y = 16'b0000001011010010;
        8: y = 16'b0000001100110100;
        9: y = 16'b0000001110010100;
        10: y = 16'b0000001111110001;
        11: y = 16'b0000010001001011;
        12: y = 16'b0000010010100011;
        13: y = 16'b0000010011110111;
        14: y = 16'b0000010101001000;
        15: y = 16'b0000010110010101;
        16: y = 16'b0000010111011111;
        17: y = 16'b0000011000100101;
        18: y = 16'b0000011001100110;
        19: y = 16'b0000011010100011;
        20: y = 16'b0000011011011100;
        21: y = 16'b0000011100010000;
        22: y = 16'b0000011100111111;
        23: y = 16'b0000011101101001;
        24: y = 16'b0000011110001110;
        25: y = 16'b0000011110101110;
        26: y = 16'b0000011111001001;
        27: y = 16'b0000011111011111;
        28: y = 16'b0000011111101111;
        29: y = 16'b0000011111111010;
        30: y = 16'b0000011111111111;
        31: y = 16'b0000011111111111;
        32: y = 16'b0000011111111010;
        33: y = 16'b0000011111101111;
        34: y = 16'b0000011111011111;
        35: y = 16'b0000011111001001;
        36: y = 16'b0000011110101110;
        37: y = 16'b0000011110001110;
        38: y = 16'b0000011101101001;
        39: y = 16'b0000011100111111;
        40: y = 16'b0000011100010000;
        41: y = 16'b0000011011011100;
        42: y = 16'b0000011010100011;
        43: y = 16'b0000011001100110;
        44: y = 16'b0000011000100101;
        45: y = 16'b0000010111011111;
        46: y = 16'b0000010110010101;
        47: y = 16'b0000010101001000;
        48: y = 16'b0000010011110111;
        49: y = 16'b0000010010100011;
        50: y = 16'b0000010001001011;
        51: y = 16'b0000001111110001;
        52: y = 16'b0000001110010100;
        53: y = 16'b0000001100110100;
        54: y = 16'b0000001011010010;
        55: y = 16'b0000001001101111;
        56: y = 16'b0000001000001010;
        57: y = 16'b0000000110100011;
        58: y = 16'b0000000100111011;
        59: y = 16'b0000000011010011;
        60: y = 16'b0000000001101001;
        61: y = 16'b0000000000000000;
        62: y = 16'b1111111110010111;
        63: y = 16'b1111111100101101;
        64: y = 16'b1111111011000101;
        65: y = 16'b1111111001011101;
        66: y = 16'b1111110111110110;
        67: y = 16'b1111110110010001;
        68: y = 16'b1111110100101110;
        69: y = 16'b1111110011001100;
        70: y = 16'b1111110001101100;
        71: y = 16'b1111110000001111;
        72: y = 16'b1111101110110101;
        73: y = 16'b1111101101011101;
        74: y = 16'b1111101100001001;
        75: y = 16'b1111101010111000;
        76: y = 16'b1111101001101011;
        77: y = 16'b1111101000100001;
        78: y = 16'b1111100111011011;
        79: y = 16'b1111100110011010;
        80: y = 16'b1111100101011101;
        81: y = 16'b1111100100100100;
        82: y = 16'b1111100011110000;
        83: y = 16'b1111100011000001;
        84: y = 16'b1111100010010111;
        85: y = 16'b1111100001110010;
        86: y = 16'b1111100001010010;
        87: y = 16'b1111100000110111;
        88: y = 16'b1111100000100001;
        89: y = 16'b1111100000010001;
        90: y = 16'b1111100000000110;
        91: y = 16'b1111100000000001;
        92: y = 16'b1111100000000001;
        93: y = 16'b1111100000000110;
        94: y = 16'b1111100000010001;
        95: y = 16'b1111100000100001;
        96: y = 16'b1111100000110111;
        97: y = 16'b1111100001010010;
        98: y = 16'b1111100001110010;
        99: y = 16'b1111100010010111;
        100: y = 16'b1111100011000001;
        101: y = 16'b1111100011110000;
        102: y = 16'b1111100100100100;
        103: y = 16'b1111100101011101;
        104: y = 16'b1111100110011010;
        105: y = 16'b1111100111011011;
        106: y = 16'b1111101000100001;
        107: y = 16'b1111101001101011;
        108: y = 16'b1111101010111000;
        109: y = 16'b1111101100001001;
        110: y = 16'b1111101101011101;
        111: y = 16'b1111101110110101;
        112: y = 16'b1111110000001111;
        113: y = 16'b1111110001101100;
        114: y = 16'b1111110011001100;
        115: y = 16'b1111110100101110;
        116: y = 16'b1111110110010001;
        117: y = 16'b1111110111110110;
        118: y = 16'b1111111001011101;
        119: y = 16'b1111111011000101;
        120: y = 16'b1111111100101101;
        121: y = 16'b1111111110010111;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=415.3Hz, Fs=48000Hz, 16-bit

module lut_Gs
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 114;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000001110000;
        2: y = 16'b0000000011011111;
        3: y = 16'b0000000101001110;
        4: y = 16'b0000000110111100;
        5: y = 16'b0000001000101001;
        6: y = 16'b0000001010010011;
        7: y = 16'b0000001011111100;
        8: y = 16'b0000001101100011;
        9: y = 16'b0000001111000111;
        10: y = 16'b0000010000101000;
        11: y = 16'b0000010010000110;
        12: y = 16'b0000010011100001;
        13: y = 16'b0000010100110111;
        14: y = 16'b0000010110001010;
        15: y = 16'b0000010111011001;
        16: y = 16'b0000011000100011;
        17: y = 16'b0000011001101000;
        18: y = 16'b0000011010101001;
        19: y = 16'b0000011011100100;
        20: y = 16'b0000011100011010;
        21: y = 16'b0000011101001011;
        22: y = 16'b0000011101110110;
        23: y = 16'b0000011110011100;
        24: y = 16'b0000011110111011;
        25: y = 16'b0000011111010101;
        26: y = 16'b0000011111101001;
        27: y = 16'b0000011111110111;
        28: y = 16'b0000011111111110;
        29: y = 16'b0000100000000000;
        30: y = 16'b0000011111111011;
        31: y = 16'b0000011111110000;
        32: y = 16'b0000011111100000;
        33: y = 16'b0000011111001001;
        34: y = 16'b0000011110101100;
        35: y = 16'b0000011110001010;
        36: y = 16'b0000011101100001;
        37: y = 16'b0000011100110011;
        38: y = 16'b0000011100000000;
        39: y = 16'b0000011011000111;
        40: y = 16'b0000011010001001;
        41: y = 16'b0000011001000110;
        42: y = 16'b0000010111111110;
        43: y = 16'b0000010110110010;
        44: y = 16'b0000010101100001;
        45: y = 16'b0000010100001100;
        46: y = 16'b0000010010110100;
        47: y = 16'b0000010001010111;
        48: y = 16'b0000001111111000;
        49: y = 16'b0000001110010101;
        50: y = 16'b0000001100110000;
        51: y = 16'b0000001011001000;
        52: y = 16'b0000001001011110;
        53: y = 16'b0000000111110010;
        54: y = 16'b0000000110000101;
        55: y = 16'b0000000100010111;
        56: y = 16'b0000000010101000;
        57: y = 16'b0000000000111000;
        58: y = 16'b1111111111001000;
        59: y = 16'b1111111101011000;
        60: y = 16'b1111111011101001;
        61: y = 16'b1111111001111011;
        62: y = 16'b1111111000001110;
        63: y = 16'b1111110110100010;
        64: y = 16'b1111110100111000;
        65: y = 16'b1111110011010000;
        66: y = 16'b1111110001101011;
        67: y = 16'b1111110000001000;
        68: y = 16'b1111101110101001;
        69: y = 16'b1111101101001100;
        70: y = 16'b1111101011110100;
        71: y = 16'b1111101010011111;
        72: y = 16'b1111101001001110;
        73: y = 16'b1111101000000010;
        74: y = 16'b1111100110111010;
        75: y = 16'b1111100101110111;
        76: y = 16'b1111100100111001;
        77: y = 16'b1111100100000000;
        78: y = 16'b1111100011001101;
        79: y = 16'b1111100010011111;
        80: y = 16'b1111100001110110;
        81: y = 16'b1111100001010100;
        82: y = 16'b1111100000110111;
        83: y = 16'b1111100000100000;
        84: y = 16'b1111100000010000;
        85: y = 16'b1111100000000101;
        86: y = 16'b1111100000000000;
        87: y = 16'b1111100000000010;
        88: y = 16'b1111100000001001;
        89: y = 16'b1111100000010111;
        90: y = 16'b1111100000101011;
        91: y = 16'b1111100001000101;
        92: y = 16'b1111100001100100;
        93: y = 16'b1111100010001010;
        94: y = 16'b1111100010110101;
        95: y = 16'b1111100011100110;
        96: y = 16'b1111100100011100;
        97: y = 16'b1111100101010111;
        98: y = 16'b1111100110011000;
        99: y = 16'b1111100111011101;
        100: y = 16'b1111101000100111;
        101: y = 16'b1111101001110110;
        102: y = 16'b1111101011001001;
        103: y = 16'b1111101100011111;
        104: y = 16'b1111101101111010;
        105: y = 16'b1111101111011000;
        106: y = 16'b1111110000111001;
        107: y = 16'b1111110010011101;
        108: y = 16'b1111110100000100;
        109: y = 16'b1111110101101101;
        110: y = 16'b1111110111010111;
        111: y = 16'b1111111001000100;
        112: y = 16'b1111111010110010;
        113: y = 16'b1111111100100001;
        114: y = 16'b1111111110010000;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=440.0Hz, Fs=48000Hz, 16-bit

module lut_A
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 108;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000001110110;
        2: y = 16'b0000000011101100;
        3: y = 16'b0000000101100000;
        4: y = 16'b0000000111010100;
        5: y = 16'b0000001001000110;
        6: y = 16'b0000001010110110;
        7: y = 16'b0000001100100100;
        8: y = 16'b0000001110001111;
        9: y = 16'b0000001111110111;
        10: y = 16'b0000010001011100;
        11: y = 16'b0000010010111101;
        12: y = 16'b0000010100011010;
        13: y = 16'b0000010101110011;
        14: y = 16'b0000010111000111;
        15: y = 16'b0000011000010110;
        16: y = 16'b0000011001100000;
        17: y = 16'b0000011010100101;
        18: y = 16'b0000011011100100;
        19: y = 16'b0000011100011101;
        20: y = 16'b0000011101010000;
        21: y = 16'b0000011101111100;
        22: y = 16'b0000011110100011;
        23: y = 16'b0000011111000011;
        24: y = 16'b0000011111011100;
        25: y = 16'b0000011111101111;
        26: y = 16'b0000011111111011;
        27: y = 16'b0000100000000000;
        28: y = 16'b0000011111111110;
        29: y = 16'b0000011111110110;
        30: y = 16'b0000011111100110;
        31: y = 16'b0000011111010000;
        32: y = 16'b0000011110110100;
        33: y = 16'b0000011110010000;
        34: y = 16'b0000011101100111;
        35: y = 16'b0000011100110111;
        36: y = 16'b0000011100000001;
        37: y = 16'b0000011011000101;
        38: y = 16'b0000011010000011;
        39: y = 16'b0000011000111100;
        40: y = 16'b0000010111101111;
        41: y = 16'b0000010110011110;
        42: y = 16'b0000010101000111;
        43: y = 16'b0000010011101100;
        44: y = 16'b0000010010001101;
        45: y = 16'b0000010000101010;
        46: y = 16'b0000001111000100;
        47: y = 16'b0000001101011010;
        48: y = 16'b0000001011101110;
        49: y = 16'b0000001001111110;
        50: y = 16'b0000001000001101;
        51: y = 16'b0000000110011010;
        52: y = 16'b0000000100100110;
        53: y = 16'b0000000010110001;
        54: y = 16'b0000000000111011;
        55: y = 16'b1111111111000101;
        56: y = 16'b1111111101001111;
        57: y = 16'b1111111011011010;
        58: y = 16'b1111111001100110;
        59: y = 16'b1111110111110011;
        60: y = 16'b1111110110000010;
        61: y = 16'b1111110100010010;
        62: y = 16'b1111110010100110;
        63: y = 16'b1111110000111100;
        64: y = 16'b1111101111010110;
        65: y = 16'b1111101101110011;
        66: y = 16'b1111101100010100;
        67: y = 16'b1111101010111001;
        68: y = 16'b1111101001100010;
        69: y = 16'b1111101000010001;
        70: y = 16'b1111100111000100;
        71: y = 16'b1111100101111101;
        72: y = 16'b1111100100111011;
        73: y = 16'b1111100011111111;
        74: y = 16'b1111100011001001;
        75: y = 16'b1111100010011001;
        76: y = 16'b1111100001110000;
        77: y = 16'b1111100001001100;
        78: y = 16'b1111100000110000;
        79: y = 16'b1111100000011010;
        80: y = 16'b1111100000001010;
        81: y = 16'b1111100000000010;
        82: y = 16'b1111100000000000;
        83: y = 16'b1111100000000101;
        84: y = 16'b1111100000010001;
        85: y = 16'b1111100000100100;
        86: y = 16'b1111100000111101;
        87: y = 16'b1111100001011101;
        88: y = 16'b1111100010000100;
        89: y = 16'b1111100010110000;
        90: y = 16'b1111100011100011;
        91: y = 16'b1111100100011100;
        92: y = 16'b1111100101011011;
        93: y = 16'b1111100110100000;
        94: y = 16'b1111100111101010;
        95: y = 16'b1111101000111001;
        96: y = 16'b1111101010001101;
        97: y = 16'b1111101011100110;
        98: y = 16'b1111101101000011;
        99: y = 16'b1111101110100100;
        100: y = 16'b1111110000001001;
        101: y = 16'b1111110001110001;
        102: y = 16'b1111110011011100;
        103: y = 16'b1111110101001010;
        104: y = 16'b1111110110111010;
        105: y = 16'b1111111000101100;
        106: y = 16'b1111111010100000;
        107: y = 16'b1111111100010100;
        108: y = 16'b1111111110001010;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=466.16Hz, Fs=48000Hz, 16-bit

module lut_As
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 101;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000001111110;
        2: y = 16'b0000000011111100;
        3: y = 16'b0000000101111000;
        4: y = 16'b0000000111110100;
        5: y = 16'b0000001001101101;
        6: y = 16'b0000001011100100;
        7: y = 16'b0000001101011000;
        8: y = 16'b0000001111001001;
        9: y = 16'b0000010000110110;
        10: y = 16'b0000010010011111;
        11: y = 16'b0000010100000100;
        12: y = 16'b0000010101100100;
        13: y = 16'b0000010110111110;
        14: y = 16'b0000011000010011;
        15: y = 16'b0000011001100010;
        16: y = 16'b0000011010101011;
        17: y = 16'b0000011011101110;
        18: y = 16'b0000011100101001;
        19: y = 16'b0000011101011110;
        20: y = 16'b0000011110001100;
        21: y = 16'b0000011110110010;
        22: y = 16'b0000011111010001;
        23: y = 16'b0000011111101000;
        24: y = 16'b0000011111110111;
        25: y = 16'b0000011111111111;
        26: y = 16'b0000011111111111;
        27: y = 16'b0000011111110111;
        28: y = 16'b0000011111101000;
        29: y = 16'b0000011111010001;
        30: y = 16'b0000011110110010;
        31: y = 16'b0000011110001100;
        32: y = 16'b0000011101011110;
        33: y = 16'b0000011100101001;
        34: y = 16'b0000011011101110;
        35: y = 16'b0000011010101011;
        36: y = 16'b0000011001100010;
        37: y = 16'b0000011000010011;
        38: y = 16'b0000010110111110;
        39: y = 16'b0000010101100100;
        40: y = 16'b0000010100000100;
        41: y = 16'b0000010010011111;
        42: y = 16'b0000010000110110;
        43: y = 16'b0000001111001001;
        44: y = 16'b0000001101011000;
        45: y = 16'b0000001011100100;
        46: y = 16'b0000001001101101;
        47: y = 16'b0000000111110100;
        48: y = 16'b0000000101111000;
        49: y = 16'b0000000011111100;
        50: y = 16'b0000000001111110;
        51: y = 16'b0000000000000000;
        52: y = 16'b1111111110000010;
        53: y = 16'b1111111100000100;
        54: y = 16'b1111111010001000;
        55: y = 16'b1111111000001100;
        56: y = 16'b1111110110010011;
        57: y = 16'b1111110100011100;
        58: y = 16'b1111110010101000;
        59: y = 16'b1111110000110111;
        60: y = 16'b1111101111001010;
        61: y = 16'b1111101101100001;
        62: y = 16'b1111101011111100;
        63: y = 16'b1111101010011100;
        64: y = 16'b1111101001000010;
        65: y = 16'b1111100111101101;
        66: y = 16'b1111100110011110;
        67: y = 16'b1111100101010101;
        68: y = 16'b1111100100010010;
        69: y = 16'b1111100011010111;
        70: y = 16'b1111100010100010;
        71: y = 16'b1111100001110100;
        72: y = 16'b1111100001001110;
        73: y = 16'b1111100000101111;
        74: y = 16'b1111100000011000;
        75: y = 16'b1111100000001001;
        76: y = 16'b1111100000000001;
        77: y = 16'b1111100000000001;
        78: y = 16'b1111100000001001;
        79: y = 16'b1111100000011000;
        80: y = 16'b1111100000101111;
        81: y = 16'b1111100001001110;
        82: y = 16'b1111100001110100;
        83: y = 16'b1111100010100010;
        84: y = 16'b1111100011010111;
        85: y = 16'b1111100100010010;
        86: y = 16'b1111100101010101;
        87: y = 16'b1111100110011110;
        88: y = 16'b1111100111101101;
        89: y = 16'b1111101001000010;
        90: y = 16'b1111101010011100;
        91: y = 16'b1111101011111100;
        92: y = 16'b1111101101100001;
        93: y = 16'b1111101111001010;
        94: y = 16'b1111110000110111;
        95: y = 16'b1111110010101000;
        96: y = 16'b1111110100011100;
        97: y = 16'b1111110110010011;
        98: y = 16'b1111111000001100;
        99: y = 16'b1111111010001000;
        100: y = 16'b1111111100000100;
        101: y = 16'b1111111110000010;
        default: y = 16'b0;
        endcase

endmodule

// y(t) = sin(2*pi*F*t), F=493.88Hz, Fs=48000Hz, 16-bit

module lut_B
(
    input        [ 7:0] x,
    output       [ 7:0] x_max,
    output logic [15:0] y
);

    assign x_max = 96;

    always_comb
        case (x)
        0: y = 16'b0000000000000000;
        1: y = 16'b0000000010000101;
        2: y = 16'b0000000100001001;
        3: y = 16'b0000000110001011;
        4: y = 16'b0000001000001101;
        5: y = 16'b0000001010001100;
        6: y = 16'b0000001100001000;
        7: y = 16'b0000001110000001;
        8: y = 16'b0000001111110110;
        9: y = 16'b0000010001100111;
        10: y = 16'b0000010011010100;
        11: y = 16'b0000010100111011;
        12: y = 16'b0000010110011100;
        13: y = 16'b0000010111111000;
        14: y = 16'b0000011001001101;
        15: y = 16'b0000011010011011;
        16: y = 16'b0000011011100010;
        17: y = 16'b0000011100100010;
        18: y = 16'b0000011101011010;
        19: y = 16'b0000011110001011;
        20: y = 16'b0000011110110011;
        21: y = 16'b0000011111010011;
        22: y = 16'b0000011111101010;
        23: y = 16'b0000011111111001;
        24: y = 16'b0000100000000000;
        25: y = 16'b0000011111111110;
        26: y = 16'b0000011111110011;
        27: y = 16'b0000011111100000;
        28: y = 16'b0000011111000100;
        29: y = 16'b0000011110100000;
        30: y = 16'b0000011101110100;
        31: y = 16'b0000011100111111;
        32: y = 16'b0000011100000011;
        33: y = 16'b0000011011000000;
        34: y = 16'b0000011001110101;
        35: y = 16'b0000011000100011;
        36: y = 16'b0000010111001011;
        37: y = 16'b0000010101101100;
        38: y = 16'b0000010100001000;
        39: y = 16'b0000010010011110;
        40: y = 16'b0000010000101111;
        41: y = 16'b0000001110111100;
        42: y = 16'b0000001101000101;
        43: y = 16'b0000001011001010;
        44: y = 16'b0000001001001101;
        45: y = 16'b0000000111001100;
        46: y = 16'b0000000101001010;
        47: y = 16'b0000000011000111;
        48: y = 16'b0000000001000010;
        49: y = 16'b1111111110111110;
        50: y = 16'b1111111100111001;
        51: y = 16'b1111111010110110;
        52: y = 16'b1111111000110100;
        53: y = 16'b1111110110110011;
        54: y = 16'b1111110100110110;
        55: y = 16'b1111110010111011;
        56: y = 16'b1111110001000100;
        57: y = 16'b1111101111010001;
        58: y = 16'b1111101101100010;
        59: y = 16'b1111101011111000;
        60: y = 16'b1111101010010100;
        61: y = 16'b1111101000110101;
        62: y = 16'b1111100111011101;
        63: y = 16'b1111100110001011;
        64: y = 16'b1111100101000000;
        65: y = 16'b1111100011111101;
        66: y = 16'b1111100011000001;
        67: y = 16'b1111100010001100;
        68: y = 16'b1111100001100000;
        69: y = 16'b1111100000111100;
        70: y = 16'b1111100000100000;
        71: y = 16'b1111100000001101;
        72: y = 16'b1111100000000010;
        73: y = 16'b1111100000000000;
        74: y = 16'b1111100000000111;
        75: y = 16'b1111100000010110;
        76: y = 16'b1111100000101101;
        77: y = 16'b1111100001001101;
        78: y = 16'b1111100001110101;
        79: y = 16'b1111100010100110;
        80: y = 16'b1111100011011110;
        81: y = 16'b1111100100011110;
        82: y = 16'b1111100101100101;
        83: y = 16'b1111100110110011;
        84: y = 16'b1111101000001000;
        85: y = 16'b1111101001100100;
        86: y = 16'b1111101011000101;
        87: y = 16'b1111101100101100;
        88: y = 16'b1111101110011001;
        89: y = 16'b1111110000001010;
        90: y = 16'b1111110001111111;
        91: y = 16'b1111110011111000;
        92: y = 16'b1111110101110100;
        93: y = 16'b1111110111110011;
        94: y = 16'b1111111001110101;
        95: y = 16'b1111111011110111;
        96: y = 16'b1111111101111011;
        default: y = 16'b0;
        endcase

endmodule

